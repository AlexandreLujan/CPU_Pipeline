library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.NUMERIC_STD.all;

entity INST_MEM is
port (
		CLOCK 	 : in  STD_LOGIC;
        ADDRESS_I: in  STD_LOGIC_VECTOR(31 downto 0);
        ADDRESS_O : out STD_LOGIC_VECTOR(31 downto 0)
     );
end INST_MEM;

architecture RTL of INST_MEM is

type rom_t is array (0 to 63) of STD_LOGIC_VECTOR(31 downto 0);
constant rom : rom_t :=
           ("01101100000000010000000000000010",  -- end 0 ADDI $A, $B, 2
            "10101100010000010000000000000000",  -- end 1 LW $C, 0($B)
            "00001000000000000000000000010000",  -- end 2 JP
            "10001100011000010000000000000000",  -- end 3 SW $D, 0($B)
            "00000000000000000000000000000000",  -- end 4
            "00000000000000000000000000000000",  -- end 5
            "00000000000000000000000000000000",  -- end 6
            "00000000000000000000000000000000",  -- end 7
            "00000000000000000000000000000000",  -- end 8
            "00000000000000000000000000000000",  -- end 9
            "00000000000000000000000000000000",  -- end 10
            "00000000000000000000000000000000",  -- end 11
            "00000000000000000000000000000000",  -- end 12
            "00000000000000000000000000000000",  -- end 13
            "00000000000000000000000000000000",  -- end 14
            "00000000000000000000000000000000",  -- end 15
            "00001100100000010000000000000110",  -- end 16
            "00000000000000000000000000000000",  -- end 17
            "00000000000000000000000000000000",  -- end 18
            "00000000000000000000000000000000",  -- end 19
            "00000000000000000000000000000000",  -- end 20
            "00000000000000000000000000000000",  -- end 21
            "00000000000000000000000000000000",  -- end 22
            "00000000000000000000000000000000",  -- end 23
            "00000000000000000000000000000000",  -- end 24
            "00000000000000000000000000000000",  -- end 25
			"00000000000000000000000000000000",  -- end 26
            "00000000000000000000000000000000",  -- end 27
            "00000000000000000000000000000000",  -- end 28
            "00000000000000000000000000000000",  -- end 29
            "00000000000000000000000000000000",  -- end 30
            "00000000000000000000000000000000",  -- end 31
			"00000000000000000000000000000000",  -- end 32
            "00000000000000000000000000000000",  -- end 33
            "00000000000000000000000000000000",  -- end 34
            "00000000000000000000000000000000",  -- end 35
            "00000000000000000000000000000000",  -- end 36
            "00000000000000000000000000000000",  -- end 37
            "00000000000000000000000000000000",  -- end 38
            "00000000000000000000000000000000",  -- end 39
            "00000000000000000000000000000000",  -- end 40
			"00000000000000000000000000000000",  -- end 41
            "00000000000000000000000000000000",  -- end 42
            "00000000000000000000000000000000",  -- end 43
            "00000000000000000000000000000000",  -- end 44
            "00000000000000000000000000000000",  -- end 45
            "00000000000000000000000000000000",  -- end 46
            "00000000000000000000000000000000",  -- end 47
            "00000000000000000000000000000000",  -- end 48
            "00000000000000000000000000000000",  -- end 49
            "00000000000000000000000000000000",  -- end 50
            "00000000000000000000000000000000",  -- end 51
			"00000000000000000000000000000000",  -- end 52
            "00000000000000000000000000000000",  -- end 53
            "00000000000000000000000000000000",  -- end 54
            "00000000000000000000000000000000",  -- end 55
            "00000000000000000000000000000000",  -- end 56
            "00000000000000000000000000000000",  -- end 57
            "00000000000000000000000000000000",  -- end 58
            "00000000000000000000000000000000",  -- end 59
            "00000000000000000000000000000000",  -- end 60
            "00000000000000000000000000000000",  -- end 61
            "00000000000000000000000000000000",  -- end 62
            "00000000000000000000000000000000"   -- end 63
);
begin

	process(CLOCK)
	begin
		if(rising_edge(CLOCK)) then
			ADDRESS_O <= rom(to_integer(signed(ADDRESS_I(31 downto 2))));
		end if;
	end process;

end RTL;
